package router_env_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
// import the YAPP package
  import yapp_pkg::*;
// other UVC packages
  import hbus_pkg::*;
  import channel_pkg::*;
  import clock_and_reset_pkg::*;	
  `include "router_reference.sv"
  `include "router_scoreboard.sv"
  `include "router_module_env.sv"  
endpackage: router_env_pkg
