// Define your enumerated type(s) here
typedef enum {GOOD_PARITY, BAD_PARITY} parity_type_e;

class yapp_packet extends uvm_sequence_item;

// Follow the lab instructions to create the packet.
// Place the packet declarations in the following order:

  // Define protocol data
  rand bit [5:0] length;
  rand bit [1:0] addr;
  rand bit [7:0] payload[];
  bit [7:0] parity;
  
  
  // Define control knobs
  rand parity_type_e parity_type;
  rand int packet_delay;
  
  // UVM_constructor for yapp_packet
  function new (string name = "yapp_packet");
    super.new(name);
  endfunction
  
  	
  // Enable automation of the packet's fields
  `uvm_object_utils_begin(yapp_packet)
  	`uvm_field_int(length,UVM_ALL_ON)
    `uvm_field_int(addr,UVM_ALL_ON)
    `uvm_field_array_int(payload,UVM_ALL_ON)
    `uvm_field_int(parity,UVM_ALL_ON)
    `uvm_field_enum(parity_type_e, parity_type, UVM_ALL_ON)
  `uvm_object_utils_end
  
  // Define packet constraints
  constraint address {addr != 3;}
  constraint payload_size {length == payload.size();}
  constraint def_length {length > 0; length < 64;}
  constraint parity_type_cons {parity_type dist {GOOD_PARITY:=8,BAD_PARITY:=2};}
  constraint packet_delay_cons {packet_delay >= 1; packet_delay <= 20;}

  // Add methods for parity calculation and class construction
  function bit [7:0] calc_parity();
    parity = {length,addr};
    
    foreach(payload[i])
      parity ^= payload[i];
    return parity;
  endfunction
  
  function void set_parity();
    if(parity_type == GOOD_PARITY)
      parity = calc_parity();
    else // if (parity_type == BAD_PARITY)
      parity = ~(calc_parity());
  endfunction
  
  function void post_randomize();
    set_parity();
  endfunction

endclass: yapp_packet


class short_yapp_packet extends yapp_packet;
  `uvm_object_utils(short_yapp_packet)
  
  function new(string name = "short_yapp_packet");
    super.new(name);
  endfunction
  
  
  
  constraint short_packet_length { length >0; length < 15;}
  //constraint address_2 { addr != 2; }
  


endclass


































